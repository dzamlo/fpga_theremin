library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity sin_lut is
port( addr: in std_logic_vector(9-1 downto 0);
      data: out signed(16-1 downto 0)
    );
end sin_lut;
architecture lut_arch of sin_lut is
begin
with addr select data <=
to_signed(0, 16) when "000000000",
to_signed(101, 16) when "000000001",
to_signed(201, 16) when "000000010",
to_signed(302, 16) when "000000011",
to_signed(403, 16) when "000000100",
to_signed(504, 16) when "000000101",
to_signed(604, 16) when "000000110",
to_signed(705, 16) when "000000111",
to_signed(806, 16) when "000001000",
to_signed(906, 16) when "000001001",
to_signed(1007, 16) when "000001010",
to_signed(1108, 16) when "000001011",
to_signed(1208, 16) when "000001100",
to_signed(1309, 16) when "000001101",
to_signed(1410, 16) when "000001110",
to_signed(1510, 16) when "000001111",
to_signed(1611, 16) when "000010000",
to_signed(1712, 16) when "000010001",
to_signed(1812, 16) when "000010010",
to_signed(1913, 16) when "000010011",
to_signed(2013, 16) when "000010100",
to_signed(2114, 16) when "000010101",
to_signed(2214, 16) when "000010110",
to_signed(2315, 16) when "000010111",
to_signed(2415, 16) when "000011000",
to_signed(2516, 16) when "000011001",
to_signed(2616, 16) when "000011010",
to_signed(2716, 16) when "000011011",
to_signed(2817, 16) when "000011100",
to_signed(2917, 16) when "000011101",
to_signed(3017, 16) when "000011110",
to_signed(3118, 16) when "000011111",
to_signed(3218, 16) when "000100000",
to_signed(3318, 16) when "000100001",
to_signed(3418, 16) when "000100010",
to_signed(3519, 16) when "000100011",
to_signed(3619, 16) when "000100100",
to_signed(3719, 16) when "000100101",
to_signed(3819, 16) when "000100110",
to_signed(3919, 16) when "000100111",
to_signed(4019, 16) when "000101000",
to_signed(4119, 16) when "000101001",
to_signed(4219, 16) when "000101010",
to_signed(4319, 16) when "000101011",
to_signed(4418, 16) when "000101100",
to_signed(4518, 16) when "000101101",
to_signed(4618, 16) when "000101110",
to_signed(4718, 16) when "000101111",
to_signed(4817, 16) when "000110000",
to_signed(4917, 16) when "000110001",
to_signed(5016, 16) when "000110010",
to_signed(5116, 16) when "000110011",
to_signed(5215, 16) when "000110100",
to_signed(5315, 16) when "000110101",
to_signed(5414, 16) when "000110110",
to_signed(5514, 16) when "000110111",
to_signed(5613, 16) when "000111000",
to_signed(5712, 16) when "000111001",
to_signed(5811, 16) when "000111010",
to_signed(5910, 16) when "000111011",
to_signed(6009, 16) when "000111100",
to_signed(6108, 16) when "000111101",
to_signed(6207, 16) when "000111110",
to_signed(6306, 16) when "000111111",
to_signed(6405, 16) when "001000000",
to_signed(6504, 16) when "001000001",
to_signed(6602, 16) when "001000010",
to_signed(6701, 16) when "001000011",
to_signed(6800, 16) when "001000100",
to_signed(6898, 16) when "001000101",
to_signed(6996, 16) when "001000110",
to_signed(7095, 16) when "001000111",
to_signed(7193, 16) when "001001000",
to_signed(7291, 16) when "001001001",
to_signed(7390, 16) when "001001010",
to_signed(7488, 16) when "001001011",
to_signed(7586, 16) when "001001100",
to_signed(7684, 16) when "001001101",
to_signed(7781, 16) when "001001110",
to_signed(7879, 16) when "001001111",
to_signed(7977, 16) when "001010000",
to_signed(8075, 16) when "001010001",
to_signed(8172, 16) when "001010010",
to_signed(8270, 16) when "001010011",
to_signed(8367, 16) when "001010100",
to_signed(8465, 16) when "001010101",
to_signed(8562, 16) when "001010110",
to_signed(8659, 16) when "001010111",
to_signed(8756, 16) when "001011000",
to_signed(8853, 16) when "001011001",
to_signed(8950, 16) when "001011010",
to_signed(9047, 16) when "001011011",
to_signed(9144, 16) when "001011100",
to_signed(9240, 16) when "001011101",
to_signed(9337, 16) when "001011110",
to_signed(9433, 16) when "001011111",
to_signed(9530, 16) when "001100000",
to_signed(9626, 16) when "001100001",
to_signed(9722, 16) when "001100010",
to_signed(9819, 16) when "001100011",
to_signed(9915, 16) when "001100100",
to_signed(10011, 16) when "001100101",
to_signed(10106, 16) when "001100110",
to_signed(10202, 16) when "001100111",
to_signed(10298, 16) when "001101000",
to_signed(10393, 16) when "001101001",
to_signed(10489, 16) when "001101010",
to_signed(10584, 16) when "001101011",
to_signed(10680, 16) when "001101100",
to_signed(10775, 16) when "001101101",
to_signed(10870, 16) when "001101110",
to_signed(10965, 16) when "001101111",
to_signed(11060, 16) when "001110000",
to_signed(11154, 16) when "001110001",
to_signed(11249, 16) when "001110010",
to_signed(11344, 16) when "001110011",
to_signed(11438, 16) when "001110100",
to_signed(11532, 16) when "001110101",
to_signed(11627, 16) when "001110110",
to_signed(11721, 16) when "001110111",
to_signed(11815, 16) when "001111000",
to_signed(11909, 16) when "001111001",
to_signed(12002, 16) when "001111010",
to_signed(12096, 16) when "001111011",
to_signed(12190, 16) when "001111100",
to_signed(12283, 16) when "001111101",
to_signed(12376, 16) when "001111110",
to_signed(12470, 16) when "001111111",
to_signed(12563, 16) when "010000000",
to_signed(12656, 16) when "010000001",
to_signed(12748, 16) when "010000010",
to_signed(12841, 16) when "010000011",
to_signed(12934, 16) when "010000100",
to_signed(13026, 16) when "010000101",
to_signed(13119, 16) when "010000110",
to_signed(13211, 16) when "010000111",
to_signed(13303, 16) when "010001000",
to_signed(13395, 16) when "010001001",
to_signed(13487, 16) when "010001010",
to_signed(13579, 16) when "010001011",
to_signed(13670, 16) when "010001100",
to_signed(13762, 16) when "010001101",
to_signed(13853, 16) when "010001110",
to_signed(13944, 16) when "010001111",
to_signed(14035, 16) when "010010000",
to_signed(14126, 16) when "010010001",
to_signed(14217, 16) when "010010010",
to_signed(14308, 16) when "010010011",
to_signed(14398, 16) when "010010100",
to_signed(14489, 16) when "010010101",
to_signed(14579, 16) when "010010110",
to_signed(14669, 16) when "010010111",
to_signed(14759, 16) when "010011000",
to_signed(14849, 16) when "010011001",
to_signed(14939, 16) when "010011010",
to_signed(15028, 16) when "010011011",
to_signed(15118, 16) when "010011100",
to_signed(15207, 16) when "010011101",
to_signed(15296, 16) when "010011110",
to_signed(15385, 16) when "010011111",
to_signed(15474, 16) when "010100000",
to_signed(15563, 16) when "010100001",
to_signed(15651, 16) when "010100010",
to_signed(15740, 16) when "010100011",
to_signed(15828, 16) when "010100100",
to_signed(15916, 16) when "010100101",
to_signed(16004, 16) when "010100110",
to_signed(16092, 16) when "010100111",
to_signed(16180, 16) when "010101000",
to_signed(16267, 16) when "010101001",
to_signed(16354, 16) when "010101010",
to_signed(16442, 16) when "010101011",
to_signed(16529, 16) when "010101100",
to_signed(16616, 16) when "010101101",
to_signed(16702, 16) when "010101110",
to_signed(16789, 16) when "010101111",
to_signed(16875, 16) when "010110000",
to_signed(16962, 16) when "010110001",
to_signed(17048, 16) when "010110010",
to_signed(17134, 16) when "010110011",
to_signed(17219, 16) when "010110100",
to_signed(17305, 16) when "010110101",
to_signed(17390, 16) when "010110110",
to_signed(17476, 16) when "010110111",
to_signed(17561, 16) when "010111000",
to_signed(17646, 16) when "010111001",
to_signed(17731, 16) when "010111010",
to_signed(17815, 16) when "010111011",
to_signed(17900, 16) when "010111100",
to_signed(17984, 16) when "010111101",
to_signed(18068, 16) when "010111110",
to_signed(18152, 16) when "010111111",
to_signed(18236, 16) when "011000000",
to_signed(18319, 16) when "011000001",
to_signed(18403, 16) when "011000010",
to_signed(18486, 16) when "011000011",
to_signed(18569, 16) when "011000100",
to_signed(18652, 16) when "011000101",
to_signed(18735, 16) when "011000110",
to_signed(18817, 16) when "011000111",
to_signed(18900, 16) when "011001000",
to_signed(18982, 16) when "011001001",
to_signed(19064, 16) when "011001010",
to_signed(19146, 16) when "011001011",
to_signed(19227, 16) when "011001100",
to_signed(19309, 16) when "011001101",
to_signed(19390, 16) when "011001110",
to_signed(19471, 16) when "011001111",
to_signed(19552, 16) when "011010000",
to_signed(19633, 16) when "011010001",
to_signed(19713, 16) when "011010010",
to_signed(19794, 16) when "011010011",
to_signed(19874, 16) when "011010100",
to_signed(19954, 16) when "011010101",
to_signed(20034, 16) when "011010110",
to_signed(20113, 16) when "011010111",
to_signed(20193, 16) when "011011000",
to_signed(20272, 16) when "011011001",
to_signed(20351, 16) when "011011010",
to_signed(20430, 16) when "011011011",
to_signed(20509, 16) when "011011100",
to_signed(20587, 16) when "011011101",
to_signed(20665, 16) when "011011110",
to_signed(20743, 16) when "011011111",
to_signed(20821, 16) when "011100000",
to_signed(20899, 16) when "011100001",
to_signed(20976, 16) when "011100010",
to_signed(21054, 16) when "011100011",
to_signed(21131, 16) when "011100100",
to_signed(21208, 16) when "011100101",
to_signed(21284, 16) when "011100110",
to_signed(21361, 16) when "011100111",
to_signed(21437, 16) when "011101000",
to_signed(21513, 16) when "011101001",
to_signed(21589, 16) when "011101010",
to_signed(21665, 16) when "011101011",
to_signed(21740, 16) when "011101100",
to_signed(21815, 16) when "011101101",
to_signed(21890, 16) when "011101110",
to_signed(21965, 16) when "011101111",
to_signed(22040, 16) when "011110000",
to_signed(22114, 16) when "011110001",
to_signed(22189, 16) when "011110010",
to_signed(22263, 16) when "011110011",
to_signed(22336, 16) when "011110100",
to_signed(22410, 16) when "011110101",
to_signed(22483, 16) when "011110110",
to_signed(22557, 16) when "011110111",
to_signed(22629, 16) when "011111000",
to_signed(22702, 16) when "011111001",
to_signed(22775, 16) when "011111010",
to_signed(22847, 16) when "011111011",
to_signed(22919, 16) when "011111100",
to_signed(22991, 16) when "011111101",
to_signed(23063, 16) when "011111110",
to_signed(23134, 16) when "011111111",
to_signed(23205, 16) when "100000000",
to_signed(23276, 16) when "100000001",
to_signed(23347, 16) when "100000010",
to_signed(23418, 16) when "100000011",
to_signed(23488, 16) when "100000100",
to_signed(23558, 16) when "100000101",
to_signed(23628, 16) when "100000110",
to_signed(23698, 16) when "100000111",
to_signed(23767, 16) when "100001000",
to_signed(23836, 16) when "100001001",
to_signed(23905, 16) when "100001010",
to_signed(23974, 16) when "100001011",
to_signed(24043, 16) when "100001100",
to_signed(24111, 16) when "100001101",
to_signed(24179, 16) when "100001110",
to_signed(24247, 16) when "100001111",
to_signed(24315, 16) when "100010000",
to_signed(24382, 16) when "100010001",
to_signed(24449, 16) when "100010010",
to_signed(24516, 16) when "100010011",
to_signed(24583, 16) when "100010100",
to_signed(24649, 16) when "100010101",
to_signed(24716, 16) when "100010110",
to_signed(24782, 16) when "100010111",
to_signed(24847, 16) when "100011000",
to_signed(24913, 16) when "100011001",
to_signed(24978, 16) when "100011010",
to_signed(25043, 16) when "100011011",
to_signed(25108, 16) when "100011100",
to_signed(25173, 16) when "100011101",
to_signed(25237, 16) when "100011110",
to_signed(25301, 16) when "100011111",
to_signed(25365, 16) when "100100000",
to_signed(25429, 16) when "100100001",
to_signed(25492, 16) when "100100010",
to_signed(25555, 16) when "100100011",
to_signed(25618, 16) when "100100100",
to_signed(25681, 16) when "100100101",
to_signed(25743, 16) when "100100110",
to_signed(25806, 16) when "100100111",
to_signed(25868, 16) when "100101000",
to_signed(25929, 16) when "100101001",
to_signed(25991, 16) when "100101010",
to_signed(26052, 16) when "100101011",
to_signed(26113, 16) when "100101100",
to_signed(26174, 16) when "100101101",
to_signed(26234, 16) when "100101110",
to_signed(26294, 16) when "100101111",
to_signed(26354, 16) when "100110000",
to_signed(26414, 16) when "100110001",
to_signed(26473, 16) when "100110010",
to_signed(26533, 16) when "100110011",
to_signed(26592, 16) when "100110100",
to_signed(26650, 16) when "100110101",
to_signed(26709, 16) when "100110110",
to_signed(26767, 16) when "100110111",
to_signed(26825, 16) when "100111000",
to_signed(26883, 16) when "100111001",
to_signed(26940, 16) when "100111010",
to_signed(26997, 16) when "100111011",
to_signed(27054, 16) when "100111100",
to_signed(27111, 16) when "100111101",
to_signed(27168, 16) when "100111110",
to_signed(27224, 16) when "100111111",
to_signed(27280, 16) when "101000000",
to_signed(27335, 16) when "101000001",
to_signed(27391, 16) when "101000010",
to_signed(27446, 16) when "101000011",
to_signed(27501, 16) when "101000100",
to_signed(27555, 16) when "101000101",
to_signed(27610, 16) when "101000110",
to_signed(27664, 16) when "101000111",
to_signed(27718, 16) when "101001000",
to_signed(27771, 16) when "101001001",
to_signed(27825, 16) when "101001010",
to_signed(27878, 16) when "101001011",
to_signed(27931, 16) when "101001100",
to_signed(27983, 16) when "101001101",
to_signed(28035, 16) when "101001110",
to_signed(28087, 16) when "101001111",
to_signed(28139, 16) when "101010000",
to_signed(28191, 16) when "101010001",
to_signed(28242, 16) when "101010010",
to_signed(28293, 16) when "101010011",
to_signed(28343, 16) when "101010100",
to_signed(28394, 16) when "101010101",
to_signed(28444, 16) when "101010110",
to_signed(28494, 16) when "101010111",
to_signed(28543, 16) when "101011000",
to_signed(28593, 16) when "101011001",
to_signed(28642, 16) when "101011010",
to_signed(28691, 16) when "101011011",
to_signed(28739, 16) when "101011100",
to_signed(28787, 16) when "101011101",
to_signed(28835, 16) when "101011110",
to_signed(28883, 16) when "101011111",
to_signed(28930, 16) when "101100000",
to_signed(28978, 16) when "101100001",
to_signed(29025, 16) when "101100010",
to_signed(29071, 16) when "101100011",
to_signed(29117, 16) when "101100100",
to_signed(29164, 16) when "101100101",
to_signed(29209, 16) when "101100110",
to_signed(29255, 16) when "101100111",
to_signed(29300, 16) when "101101000",
to_signed(29345, 16) when "101101001",
to_signed(29390, 16) when "101101010",
to_signed(29434, 16) when "101101011",
to_signed(29478, 16) when "101101100",
to_signed(29522, 16) when "101101101",
to_signed(29566, 16) when "101101110",
to_signed(29609, 16) when "101101111",
to_signed(29652, 16) when "101110000",
to_signed(29695, 16) when "101110001",
to_signed(29737, 16) when "101110010",
to_signed(29779, 16) when "101110011",
to_signed(29821, 16) when "101110100",
to_signed(29863, 16) when "101110101",
to_signed(29904, 16) when "101110110",
to_signed(29945, 16) when "101110111",
to_signed(29986, 16) when "101111000",
to_signed(30026, 16) when "101111001",
to_signed(30066, 16) when "101111010",
to_signed(30106, 16) when "101111011",
to_signed(30146, 16) when "101111100",
to_signed(30185, 16) when "101111101",
to_signed(30224, 16) when "101111110",
to_signed(30263, 16) when "101111111",
to_signed(30302, 16) when "110000000",
to_signed(30340, 16) when "110000001",
to_signed(30378, 16) when "110000010",
to_signed(30415, 16) when "110000011",
to_signed(30453, 16) when "110000100",
to_signed(30490, 16) when "110000101",
to_signed(30526, 16) when "110000110",
to_signed(30563, 16) when "110000111",
to_signed(30599, 16) when "110001000",
to_signed(30635, 16) when "110001001",
to_signed(30671, 16) when "110001010",
to_signed(30706, 16) when "110001011",
to_signed(30741, 16) when "110001100",
to_signed(30776, 16) when "110001101",
to_signed(30810, 16) when "110001110",
to_signed(30844, 16) when "110001111",
to_signed(30878, 16) when "110010000",
to_signed(30912, 16) when "110010001",
to_signed(30945, 16) when "110010010",
to_signed(30978, 16) when "110010011",
to_signed(31010, 16) when "110010100",
to_signed(31043, 16) when "110010101",
to_signed(31075, 16) when "110010110",
to_signed(31107, 16) when "110010111",
to_signed(31138, 16) when "110011000",
to_signed(31169, 16) when "110011001",
to_signed(31200, 16) when "110011010",
to_signed(31231, 16) when "110011011",
to_signed(31261, 16) when "110011100",
to_signed(31291, 16) when "110011101",
to_signed(31321, 16) when "110011110",
to_signed(31351, 16) when "110011111",
to_signed(31380, 16) when "110100000",
to_signed(31409, 16) when "110100001",
to_signed(31437, 16) when "110100010",
to_signed(31465, 16) when "110100011",
to_signed(31493, 16) when "110100100",
to_signed(31521, 16) when "110100101",
to_signed(31548, 16) when "110100110",
to_signed(31575, 16) when "110100111",
to_signed(31602, 16) when "110101000",
to_signed(31629, 16) when "110101001",
to_signed(31655, 16) when "110101010",
to_signed(31681, 16) when "110101011",
to_signed(31706, 16) when "110101100",
to_signed(31732, 16) when "110101101",
to_signed(31757, 16) when "110101110",
to_signed(31781, 16) when "110101111",
to_signed(31806, 16) when "110110000",
to_signed(31830, 16) when "110110001",
to_signed(31853, 16) when "110110010",
to_signed(31877, 16) when "110110011",
to_signed(31900, 16) when "110110100",
to_signed(31923, 16) when "110110101",
to_signed(31945, 16) when "110110110",
to_signed(31968, 16) when "110110111",
to_signed(31990, 16) when "110111000",
to_signed(32011, 16) when "110111001",
to_signed(32033, 16) when "110111010",
to_signed(32054, 16) when "110111011",
to_signed(32075, 16) when "110111100",
to_signed(32095, 16) when "110111101",
to_signed(32115, 16) when "110111110",
to_signed(32135, 16) when "110111111",
to_signed(32154, 16) when "111000000",
to_signed(32174, 16) when "111000001",
to_signed(32193, 16) when "111000010",
to_signed(32211, 16) when "111000011",
to_signed(32230, 16) when "111000100",
to_signed(32248, 16) when "111000101",
to_signed(32265, 16) when "111000110",
to_signed(32283, 16) when "111000111",
to_signed(32300, 16) when "111001000",
to_signed(32317, 16) when "111001001",
to_signed(32333, 16) when "111001010",
to_signed(32349, 16) when "111001011",
to_signed(32365, 16) when "111001100",
to_signed(32381, 16) when "111001101",
to_signed(32396, 16) when "111001110",
to_signed(32411, 16) when "111001111",
to_signed(32426, 16) when "111010000",
to_signed(32440, 16) when "111010001",
to_signed(32454, 16) when "111010010",
to_signed(32468, 16) when "111010011",
to_signed(32481, 16) when "111010100",
to_signed(32494, 16) when "111010101",
to_signed(32507, 16) when "111010110",
to_signed(32520, 16) when "111010111",
to_signed(32532, 16) when "111011000",
to_signed(32544, 16) when "111011001",
to_signed(32555, 16) when "111011010",
to_signed(32567, 16) when "111011011",
to_signed(32578, 16) when "111011100",
to_signed(32588, 16) when "111011101",
to_signed(32599, 16) when "111011110",
to_signed(32609, 16) when "111011111",
to_signed(32618, 16) when "111100000",
to_signed(32628, 16) when "111100001",
to_signed(32637, 16) when "111100010",
to_signed(32646, 16) when "111100011",
to_signed(32654, 16) when "111100100",
to_signed(32662, 16) when "111100101",
to_signed(32670, 16) when "111100110",
to_signed(32678, 16) when "111100111",
to_signed(32685, 16) when "111101000",
to_signed(32692, 16) when "111101001",
to_signed(32699, 16) when "111101010",
to_signed(32705, 16) when "111101011",
to_signed(32711, 16) when "111101100",
to_signed(32717, 16) when "111101101",
to_signed(32722, 16) when "111101110",
to_signed(32727, 16) when "111101111",
to_signed(32732, 16) when "111110000",
to_signed(32737, 16) when "111110001",
to_signed(32741, 16) when "111110010",
to_signed(32745, 16) when "111110011",
to_signed(32748, 16) when "111110100",
to_signed(32752, 16) when "111110101",
to_signed(32754, 16) when "111110110",
to_signed(32757, 16) when "111110111",
to_signed(32759, 16) when "111111000",
to_signed(32761, 16) when "111111001",
to_signed(32763, 16) when "111111010",
to_signed(32765, 16) when "111111011",
to_signed(32766, 16) when "111111100",
to_signed(32766, 16) when "111111101",
to_signed(32767, 16) when "111111110",
to_signed(32767, 16) when "111111111",
to_signed(0, 16) when others;
end lut_arch;

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity dist_correct is
port( addr: in std_logic_vector(8-1 downto 0);
      data: out unsigned(8-1 downto 0)
    );
end dist_correct;
architecture lut_arch of dist_correct is
begin
with addr select data <=
to_unsigned(0, 8) when "00000000",
to_unsigned(1, 8) when "00000001",
to_unsigned(3, 8) when "00000010",
to_unsigned(4, 8) when "00000011",
to_unsigned(5, 8) when "00000100",
to_unsigned(7, 8) when "00000101",
to_unsigned(8, 8) when "00000110",
to_unsigned(9, 8) when "00000111",
to_unsigned(11, 8) when "00001000",
to_unsigned(12, 8) when "00001001",
to_unsigned(13, 8) when "00001010",
to_unsigned(15, 8) when "00001011",
to_unsigned(16, 8) when "00001100",
to_unsigned(17, 8) when "00001101",
to_unsigned(18, 8) when "00001110",
to_unsigned(20, 8) when "00001111",
to_unsigned(21, 8) when "00010000",
to_unsigned(22, 8) when "00010001",
to_unsigned(24, 8) when "00010010",
to_unsigned(25, 8) when "00010011",
to_unsigned(26, 8) when "00010100",
to_unsigned(28, 8) when "00010101",
to_unsigned(29, 8) when "00010110",
to_unsigned(30, 8) when "00010111",
to_unsigned(32, 8) when "00011000",
to_unsigned(33, 8) when "00011001",
to_unsigned(34, 8) when "00011010",
to_unsigned(36, 8) when "00011011",
to_unsigned(37, 8) when "00011100",
to_unsigned(38, 8) when "00011101",
to_unsigned(40, 8) when "00011110",
to_unsigned(41, 8) when "00011111",
to_unsigned(42, 8) when "00100000",
to_unsigned(44, 8) when "00100001",
to_unsigned(45, 8) when "00100010",
to_unsigned(46, 8) when "00100011",
to_unsigned(48, 8) when "00100100",
to_unsigned(49, 8) when "00100101",
to_unsigned(50, 8) when "00100110",
to_unsigned(52, 8) when "00100111",
to_unsigned(53, 8) when "00101000",
to_unsigned(54, 8) when "00101001",
to_unsigned(55, 8) when "00101010",
to_unsigned(57, 8) when "00101011",
to_unsigned(58, 8) when "00101100",
to_unsigned(59, 8) when "00101101",
to_unsigned(61, 8) when "00101110",
to_unsigned(62, 8) when "00101111",
to_unsigned(63, 8) when "00110000",
to_unsigned(65, 8) when "00110001",
to_unsigned(66, 8) when "00110010",
to_unsigned(67, 8) when "00110011",
to_unsigned(69, 8) when "00110100",
to_unsigned(70, 8) when "00110101",
to_unsigned(71, 8) when "00110110",
to_unsigned(73, 8) when "00110111",
to_unsigned(74, 8) when "00111000",
to_unsigned(75, 8) when "00111001",
to_unsigned(77, 8) when "00111010",
to_unsigned(78, 8) when "00111011",
to_unsigned(79, 8) when "00111100",
to_unsigned(81, 8) when "00111101",
to_unsigned(82, 8) when "00111110",
to_unsigned(83, 8) when "00111111",
to_unsigned(85, 8) when "01000000",
to_unsigned(86, 8) when "01000001",
to_unsigned(87, 8) when "01000010",
to_unsigned(89, 8) when "01000011",
to_unsigned(90, 8) when "01000100",
to_unsigned(91, 8) when "01000101",
to_unsigned(92, 8) when "01000110",
to_unsigned(94, 8) when "01000111",
to_unsigned(95, 8) when "01001000",
to_unsigned(96, 8) when "01001001",
to_unsigned(98, 8) when "01001010",
to_unsigned(99, 8) when "01001011",
to_unsigned(100, 8) when "01001100",
to_unsigned(102, 8) when "01001101",
to_unsigned(103, 8) when "01001110",
to_unsigned(104, 8) when "01001111",
to_unsigned(106, 8) when "01010000",
to_unsigned(107, 8) when "01010001",
to_unsigned(108, 8) when "01010010",
to_unsigned(110, 8) when "01010011",
to_unsigned(111, 8) when "01010100",
to_unsigned(112, 8) when "01010101",
to_unsigned(114, 8) when "01010110",
to_unsigned(115, 8) when "01010111",
to_unsigned(116, 8) when "01011000",
to_unsigned(118, 8) when "01011001",
to_unsigned(119, 8) when "01011010",
to_unsigned(120, 8) when "01011011",
to_unsigned(122, 8) when "01011100",
to_unsigned(123, 8) when "01011101",
to_unsigned(124, 8) when "01011110",
to_unsigned(126, 8) when "01011111",
to_unsigned(127, 8) when "01100000",
to_unsigned(128, 8) when "01100001",
to_unsigned(129, 8) when "01100010",
to_unsigned(131, 8) when "01100011",
to_unsigned(132, 8) when "01100100",
to_unsigned(133, 8) when "01100101",
to_unsigned(135, 8) when "01100110",
to_unsigned(136, 8) when "01100111",
to_unsigned(137, 8) when "01101000",
to_unsigned(139, 8) when "01101001",
to_unsigned(140, 8) when "01101010",
to_unsigned(141, 8) when "01101011",
to_unsigned(143, 8) when "01101100",
to_unsigned(144, 8) when "01101101",
to_unsigned(145, 8) when "01101110",
to_unsigned(147, 8) when "01101111",
to_unsigned(148, 8) when "01110000",
to_unsigned(149, 8) when "01110001",
to_unsigned(151, 8) when "01110010",
to_unsigned(152, 8) when "01110011",
to_unsigned(153, 8) when "01110100",
to_unsigned(155, 8) when "01110101",
to_unsigned(156, 8) when "01110110",
to_unsigned(157, 8) when "01110111",
to_unsigned(159, 8) when "01111000",
to_unsigned(160, 8) when "01111001",
to_unsigned(161, 8) when "01111010",
to_unsigned(163, 8) when "01111011",
to_unsigned(164, 8) when "01111100",
to_unsigned(165, 8) when "01111101",
to_unsigned(166, 8) when "01111110",
to_unsigned(168, 8) when "01111111",
to_unsigned(169, 8) when "10000000",
to_unsigned(170, 8) when "10000001",
to_unsigned(172, 8) when "10000010",
to_unsigned(173, 8) when "10000011",
to_unsigned(174, 8) when "10000100",
to_unsigned(176, 8) when "10000101",
to_unsigned(177, 8) when "10000110",
to_unsigned(178, 8) when "10000111",
to_unsigned(180, 8) when "10001000",
to_unsigned(181, 8) when "10001001",
to_unsigned(182, 8) when "10001010",
to_unsigned(184, 8) when "10001011",
to_unsigned(185, 8) when "10001100",
to_unsigned(186, 8) when "10001101",
to_unsigned(188, 8) when "10001110",
to_unsigned(189, 8) when "10001111",
to_unsigned(190, 8) when "10010000",
to_unsigned(192, 8) when "10010001",
to_unsigned(193, 8) when "10010010",
to_unsigned(194, 8) when "10010011",
to_unsigned(196, 8) when "10010100",
to_unsigned(197, 8) when "10010101",
to_unsigned(198, 8) when "10010110",
to_unsigned(200, 8) when "10010111",
to_unsigned(201, 8) when "10011000",
to_unsigned(202, 8) when "10011001",
to_unsigned(203, 8) when "10011010",
to_unsigned(205, 8) when "10011011",
to_unsigned(206, 8) when "10011100",
to_unsigned(207, 8) when "10011101",
to_unsigned(209, 8) when "10011110",
to_unsigned(210, 8) when "10011111",
to_unsigned(211, 8) when "10100000",
to_unsigned(213, 8) when "10100001",
to_unsigned(214, 8) when "10100010",
to_unsigned(215, 8) when "10100011",
to_unsigned(217, 8) when "10100100",
to_unsigned(218, 8) when "10100101",
to_unsigned(219, 8) when "10100110",
to_unsigned(221, 8) when "10100111",
to_unsigned(222, 8) when "10101000",
to_unsigned(223, 8) when "10101001",
to_unsigned(225, 8) when "10101010",
to_unsigned(226, 8) when "10101011",
to_unsigned(227, 8) when "10101100",
to_unsigned(229, 8) when "10101101",
to_unsigned(230, 8) when "10101110",
to_unsigned(231, 8) when "10101111",
to_unsigned(233, 8) when "10110000",
to_unsigned(234, 8) when "10110001",
to_unsigned(235, 8) when "10110010",
to_unsigned(237, 8) when "10110011",
to_unsigned(238, 8) when "10110100",
to_unsigned(239, 8) when "10110101",
to_unsigned(240, 8) when "10110110",
to_unsigned(242, 8) when "10110111",
to_unsigned(243, 8) when "10111000",
to_unsigned(244, 8) when "10111001",
to_unsigned(246, 8) when "10111010",
to_unsigned(247, 8) when "10111011",
to_unsigned(248, 8) when "10111100",
to_unsigned(250, 8) when "10111101",
to_unsigned(251, 8) when "10111110",
to_unsigned(252, 8) when "10111111",
to_unsigned(254, 8) when "11000000",
to_unsigned(255, 8) when "11000001",
to_unsigned(256, 8) when "11000010",
to_unsigned(258, 8) when "11000011",
to_unsigned(259, 8) when "11000100",
to_unsigned(260, 8) when "11000101",
to_unsigned(262, 8) when "11000110",
to_unsigned(263, 8) when "11000111",
to_unsigned(264, 8) when "11001000",
to_unsigned(266, 8) when "11001001",
to_unsigned(267, 8) when "11001010",
to_unsigned(268, 8) when "11001011",
to_unsigned(270, 8) when "11001100",
to_unsigned(271, 8) when "11001101",
to_unsigned(272, 8) when "11001110",
to_unsigned(273, 8) when "11001111",
to_unsigned(275, 8) when "11010000",
to_unsigned(276, 8) when "11010001",
to_unsigned(277, 8) when "11010010",
to_unsigned(279, 8) when "11010011",
to_unsigned(280, 8) when "11010100",
to_unsigned(281, 8) when "11010101",
to_unsigned(283, 8) when "11010110",
to_unsigned(284, 8) when "11010111",
to_unsigned(285, 8) when "11011000",
to_unsigned(287, 8) when "11011001",
to_unsigned(288, 8) when "11011010",
to_unsigned(289, 8) when "11011011",
to_unsigned(291, 8) when "11011100",
to_unsigned(292, 8) when "11011101",
to_unsigned(293, 8) when "11011110",
to_unsigned(295, 8) when "11011111",
to_unsigned(296, 8) when "11100000",
to_unsigned(297, 8) when "11100001",
to_unsigned(299, 8) when "11100010",
to_unsigned(300, 8) when "11100011",
to_unsigned(301, 8) when "11100100",
to_unsigned(303, 8) when "11100101",
to_unsigned(304, 8) when "11100110",
to_unsigned(305, 8) when "11100111",
to_unsigned(307, 8) when "11101000",
to_unsigned(308, 8) when "11101001",
to_unsigned(309, 8) when "11101010",
to_unsigned(310, 8) when "11101011",
to_unsigned(312, 8) when "11101100",
to_unsigned(313, 8) when "11101101",
to_unsigned(314, 8) when "11101110",
to_unsigned(316, 8) when "11101111",
to_unsigned(317, 8) when "11110000",
to_unsigned(318, 8) when "11110001",
to_unsigned(320, 8) when "11110010",
to_unsigned(321, 8) when "11110011",
to_unsigned(322, 8) when "11110100",
to_unsigned(324, 8) when "11110101",
to_unsigned(325, 8) when "11110110",
to_unsigned(326, 8) when "11110111",
to_unsigned(328, 8) when "11111000",
to_unsigned(329, 8) when "11111001",
to_unsigned(330, 8) when "11111010",
to_unsigned(332, 8) when "11111011",
to_unsigned(333, 8) when "11111100",
to_unsigned(334, 8) when "11111101",
to_unsigned(336, 8) when "11111110",
to_unsigned(337, 8) when "11111111",
to_unsigned(0, 8) when others;
end lut_arch;
